module fp_mul_checker (
    input logic [31:0] fp_X,
    input logic [31:0] fp_Y,
    input logic [31:0] fp_Z,
    input logic [2:0] r_mode,
    input logic       ovrf, 
    input logic       udrf
);
endmodule
bind fp_adder fp_adder_checker chk (
  .fp_a(fp_a),
  .fp_b(fp_b),
  .r_mode(r_mode),
  .fp_result(fp_result),
  .overflow(overflow),
  .underflow(underflow)
);

// Bind del assertions al DUT
bind fp_alu alu_assertions checker_inst (.*);
